* SPICE модель выходной цепи микропередатчика

* источник питания +3.3В (пока не используется)
* VCC vcc 0 DC 3.3V

* источник синусоидального сигнала (амплитуда = 1В)
VSIN vin 0 dc 0 ac 1V sin(0 1V 433MegHz)

* сопротивление источника
R0 vin v0 10

* нагрузка (активное сопротивление "элекрростатической" антенны)
RA vout 0 10k

* индуктивности
L1 0   v0   56n
L2 v1  v2   12n
L3 v2  0    12n
L4 v3  vout 127n

* конденсаторы
C1 v0   v1 100p
C2 v2   0  10p
C3 v2   v3 33p
C4 v3   0  16p
C5 vout 0  1p

* температурный режим
.options TEMP=25

* моделирование переходного процесса
* шаг моделирования - 5 пс
* время моделирования - 30 нс
.tran 5p 30n

.end




